//    Modifications made by Praveen S G in 2024.

// Copyright 2023 MERL-DSU

//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at

//        http://www.apache.org/licenses/LICENSE-2.0

//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.

module Instruction_Memory(rst, A, RD);

  // Inputs
  input rst;                        // Reset signal
  input [31:0] A;                   // Instruction address

  // Output
  output [31:0] RD;                 // Instruction data output

  reg [31:0] mem [1023:0];          // Memory array (1K x 32-bit)

  // Read instruction from memory
  // If reset is low, output zero, otherwise read from memory
  assign RD = (rst == 1'b0) ? {32{1'b0}} : mem[A[31:2]];

  // Initialize memory contents from a hex file (memfile.hex)
  initial begin
    $readmemh("memfile.hex", mem);
  end

/*
  Example manual initialization of memory (commented out)
  initial begin
    // mem[0] = 32'hFFC4A303;
    // mem[1] = 32'h00832383;
    mem[0] = 32'h0062E233;
    // mem[1] = 32'h00B62423;
  end
*/

endmodule
